`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:04:21 11/21/2018 
// Design Name: 
// Module Name:    CodeMem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CodeMem(
    input [31:0] pc,
    output [31:0] instr
    );
	reg[31:0] code_mem[0:255];
	
	reg[31:0] instr_reg;
	assign instr = instr_reg;
	
	always@(pc)
		instr_reg = code_mem[pc];
		
    initial
        begin
            code_mem[0] <= 32'b00000000000000000000000000000010;
            code_mem[1] <= 32'b00000100001000000001000000000000;
            code_mem[2] <= 32'b00000100001000000001000000000000;
            code_mem[3] <= 32'b00001000001000100001100000000000;
            code_mem[4] <= 32'b00010100001000010000000000000000;
            code_mem[5] <= 32'b00001100011000010000000000000000;
            code_mem[6] <= 32'b00010000001000100000000000000000;
            code_mem[7] <= 32'b00011000001001000010100000000000;
            code_mem[8] <= 32'b00000101010000000000000000000000;
            code_mem[9] <= 32'b10000100000000000000000000000010;
            code_mem[10] <= 32'b00000101011000000000000000000000;
            code_mem[11] <= 32'b00100100001000000000000000000000;
            code_mem[12] <= 32'b00000101011000000000000000000000;
            code_mem[13] <= 32'b00100100001000000000000000000000;
            code_mem[14] <= 32'b01000101100000000000000000000000;
            code_mem[15] <= 32'b00000000000000000000000000000000;
            code_mem[16] <= 32'b00000000000000000000000000000000;
            code_mem[17] <= 32'b00000000000000000000000000000000;
            code_mem[18] <= 32'b00000000000000000000000000000000;
            code_mem[19] <= 32'b00000000000000000000000000000000;
            code_mem[20] <= 32'b00000000000000000000000000000000;
            code_mem[21] <= 32'b00000000000000000000000000000000;
            code_mem[22] <= 32'b00000000000000000000000000000000;
            code_mem[23] <= 32'b00000000000000000000000000000000;
            code_mem[24] <= 32'b00000000000000000000000000000000;
            code_mem[25] <= 32'b00000000000000000000000000000000;
            code_mem[26] <= 32'b00000000000000000000000000000000;
            code_mem[27] <= 32'b00000000000000000000000000000000;
            code_mem[28] <= 32'b00000000000000000000000000000000;
            code_mem[29] <= 32'b00000000000000000000000000000000;
            code_mem[30] <= 32'b00000000000000000000000000000000;
            code_mem[31] <= 32'b00000000000000000000000000000000;
            code_mem[32] <= 32'b00000000000000000000000000000000;
            code_mem[33] <= 32'b00000000000000000000000000000000;
            code_mem[34] <= 32'b00000000000000000000000000000000;
            code_mem[35] <= 32'b00000000000000000000000000000000;
            code_mem[36] <= 32'b00000000000000000000000000000000;
            code_mem[37] <= 32'b00000000000000000000000000000000;
            code_mem[38] <= 32'b00000000000000000000000000000000;
            code_mem[39] <= 32'b00000000000000000000000000000000;
            code_mem[40] <= 32'b00000000000000000000000000000000;
            code_mem[41] <= 32'b00000000000000000000000000000000;
            code_mem[42] <= 32'b00000000000000000000000000000000;
            code_mem[43] <= 32'b00000000000000000000000000000000;
            code_mem[44] <= 32'b00000000000000000000000000000000;
            code_mem[45] <= 32'b00000000000000000000000000000000;
            code_mem[46] <= 32'b00000000000000000000000000000000;
            code_mem[47] <= 32'b00000000000000000000000000000000;
            code_mem[48] <= 32'b00000000000000000000000000000000;
            code_mem[49] <= 32'b00000000000000000000000000000000;
            code_mem[50] <= 32'b00000000000000000000000000000000;
            code_mem[51] <= 32'b00000000000000000000000000000000;
            code_mem[52] <= 32'b00000000000000000000000000000000;
            code_mem[53] <= 32'b00000000000000000000000000000000;
            code_mem[54] <= 32'b00000000000000000000000000000000;
            code_mem[55] <= 32'b00000000000000000000000000000000;
            code_mem[56] <= 32'b00000000000000000000000000000000;
            code_mem[57] <= 32'b00000000000000000000000000000000;
            code_mem[58] <= 32'b00000000000000000000000000000000;
            code_mem[59] <= 32'b00000000000000000000000000000000;
            code_mem[60] <= 32'b00000000000000000000000000000000;
            code_mem[61] <= 32'b00000000000000000000000000000000;
            code_mem[62] <= 32'b00000000000000000000000000000000;
            code_mem[63] <= 32'b00000000000000000000000000000000;
            code_mem[64] <= 32'b00000000000000000000000000000000;
            code_mem[65] <= 32'b00000000000000000000000000000000;
            code_mem[66] <= 32'b00000000000000000000000000000000;
            code_mem[67] <= 32'b00000000000000000000000000000000;
            code_mem[68] <= 32'b00000000000000000000000000000000;
            code_mem[69] <= 32'b00000000000000000000000000000000;
            code_mem[70] <= 32'b00000000000000000000000000000000;
            code_mem[71] <= 32'b00000000000000000000000000000000;
            code_mem[72] <= 32'b00000000000000000000000000000000;
            code_mem[73] <= 32'b00000000000000000000000000000000;
            code_mem[74] <= 32'b00000000000000000000000000000000;
            code_mem[75] <= 32'b00000000000000000000000000000000;
            code_mem[76] <= 32'b00000000000000000000000000000000;
            code_mem[77] <= 32'b00000000000000000000000000000000;
            code_mem[78] <= 32'b00000000000000000000000000000000;
            code_mem[79] <= 32'b00000000000000000000000000000000;
            code_mem[80] <= 32'b00000000000000000000000000000000;
            code_mem[81] <= 32'b00000000000000000000000000000000;
            code_mem[82] <= 32'b00000000000000000000000000000000;
            code_mem[83] <= 32'b00000000000000000000000000000000;
            code_mem[84] <= 32'b00000000000000000000000000000000;
            code_mem[85] <= 32'b00000000000000000000000000000000;
            code_mem[86] <= 32'b00000000000000000000000000000000;
            code_mem[87] <= 32'b00000000000000000000000000000000;
            code_mem[88] <= 32'b00000000000000000000000000000000;
            code_mem[89] <= 32'b00000000000000000000000000000000;
            code_mem[90] <= 32'b00000000000000000000000000000000;
            code_mem[91] <= 32'b00000000000000000000000000000000;
            code_mem[92] <= 32'b00000000000000000000000000000000;
            code_mem[93] <= 32'b00000000000000000000000000000000;
            code_mem[94] <= 32'b00000000000000000000000000000000;
            code_mem[95] <= 32'b00000000000000000000000000000000;
            code_mem[96] <= 32'b00000000000000000000000000000000;
            code_mem[97] <= 32'b00000000000000000000000000000000;
            code_mem[98] <= 32'b00000000000000000000000000000000;
            code_mem[99] <= 32'b00000000000000000000000000000000;
            code_mem[100] <= 32'b00000000000000000000000000000000;
            code_mem[101] <= 32'b00000000000000000000000000000000;
            code_mem[102] <= 32'b00000000000000000000000000000000;
            code_mem[103] <= 32'b00000000000000000000000000000000;
            code_mem[104] <= 32'b00000000000000000000000000000000;
            code_mem[105] <= 32'b00000000000000000000000000000000;
            code_mem[106] <= 32'b00000000000000000000000000000000;
            code_mem[107] <= 32'b00000000000000000000000000000000;
            code_mem[108] <= 32'b00000000000000000000000000000000;
            code_mem[109] <= 32'b00000000000000000000000000000000;
            code_mem[110] <= 32'b00000000000000000000000000000000;
            code_mem[111] <= 32'b00000000000000000000000000000000;
            code_mem[112] <= 32'b00000000000000000000000000000000;
            code_mem[113] <= 32'b00000000000000000000000000000000;
            code_mem[114] <= 32'b00000000000000000000000000000000;
            code_mem[115] <= 32'b00000000000000000000000000000000;
            code_mem[116] <= 32'b00000000000000000000000000000000;
            code_mem[117] <= 32'b00000000000000000000000000000000;
            code_mem[118] <= 32'b00000000000000000000000000000000;
            code_mem[119] <= 32'b00000000000000000000000000000000;
            code_mem[120] <= 32'b00000000000000000000000000000000;
            code_mem[121] <= 32'b00000000000000000000000000000000;
            code_mem[122] <= 32'b00000000000000000000000000000000;
            code_mem[123] <= 32'b00000000000000000000000000000000;
            code_mem[124] <= 32'b00000000000000000000000000000000;
            code_mem[125] <= 32'b00000000000000000000000000000000;
            code_mem[126] <= 32'b00000000000000000000000000000000;
            code_mem[127] <= 32'b00000000000000000000000000000000;
            code_mem[128] <= 32'b00000000000000000000000000000000;
            code_mem[129] <= 32'b00000100001000000000000000000000;
            code_mem[130] <= 32'b00000100010000000000000000000000;
            code_mem[131] <= 32'b00010100011000000000000000000000;
            code_mem[132] <= 32'b00011000010000000001100000000000;
            code_mem[133] <= 32'b00000100011000000001000000000000;
            code_mem[134] <= 32'b00000100010000100001000000000000;
            code_mem[135] <= 32'b00000100010000100001000000000000;
            code_mem[136] <= 32'b00000100010000100001000000000000;
            code_mem[137] <= 32'b00000100010000100001000000000000;
            code_mem[138] <= 32'b00000100010000100001000000000000;
            code_mem[139] <= 32'b00000100010000100001000000000000;
            code_mem[140] <= 32'b00000100010000100001000000000000;
            code_mem[141] <= 32'b00000100010000100001000000000000;
            code_mem[142] <= 32'b00100100000000010000000000000000;
            code_mem[143] <= 32'b00000100001000010001100000000000;
            code_mem[144] <= 32'b10000100001000100000000000000010;
            code_mem[145] <= 32'b00000000000000000000000010001101;
            code_mem[146] <= 32'b00000100001000000000000000000000;
            code_mem[147] <= 32'b00000100010000000000000000000000;
            code_mem[148] <= 32'b00000100011000000000000000000000;
            code_mem[149] <= 32'b00000100100000000000000000000000;
            code_mem[150] <= 32'b00000100101000000000000000000000;
            code_mem[151] <= 32'b00000100110000000000000000000000;
            code_mem[152] <= 32'b00000100111000000000000000000000;
            code_mem[153] <= 32'b00000101000000000000000000000000;
            code_mem[154] <= 32'b00000101001000000000000000000000;
            code_mem[155] <= 32'b00000101010000000000000000000000;
            code_mem[156] <= 32'b00000101011000000000000000000000;
            code_mem[157] <= 32'b00000101100000000000000000000000;
            code_mem[158] <= 32'b00000101101000000000000000000000;
            code_mem[159] <= 32'b00000101110000000000000000000000;
            code_mem[160] <= 32'b00000101111000000000000000000000;
            code_mem[161] <= 32'b00000110000000000000000000000000;
            code_mem[162] <= 32'b00000110001000000000000000000000;
            code_mem[163] <= 32'b00000110010000000000000000000000;
            code_mem[164] <= 32'b00000110011000000000000000000000;
            code_mem[165] <= 32'b00000110100000000000000000000000;
            code_mem[166] <= 32'b00000110101000000000000000000000;
            code_mem[167] <= 32'b00000110110000000000000000000000;
            code_mem[168] <= 32'b00000110111000000000000000000000;
            code_mem[169] <= 32'b00000111000000000000000000000000;
            code_mem[170] <= 32'b00000111001000000000000000000000;
            code_mem[171] <= 32'b00000111010000000000000000000000;
            code_mem[172] <= 32'b00000111011000000000000000000000;
            code_mem[173] <= 32'b00000111100000000000000000000000;
            code_mem[174] <= 32'b00000111101000000000000000000000;
            code_mem[175] <= 32'b00000111110000000000000000000000;
            code_mem[176] <= 32'b00000111111000000000000000000000;
            code_mem[177] <= 32'b00000000000000000000000000000000;
            code_mem[178] <= 32'b00000000000000000000000000000000;
            code_mem[179] <= 32'b00000000000000000000000000000000;
            code_mem[180] <= 32'b00000000000000000000000000000000;
            code_mem[181] <= 32'b00000000000000000000000000000000;
            code_mem[182] <= 32'b00000000000000000000000000000000;
            code_mem[183] <= 32'b00000000000000000000000000000000;
            code_mem[184] <= 32'b00000000000000000000000000000000;
            code_mem[185] <= 32'b00000000000000000000000000000000;
            code_mem[186] <= 32'b00000000000000000000000000000000;
            code_mem[187] <= 32'b00000000000000000000000000000000;
            code_mem[188] <= 32'b00000000000000000000000000000000;
            code_mem[189] <= 32'b00000000000000000000000000000000;
            code_mem[190] <= 32'b00000000000000000000000000000000;
            code_mem[191] <= 32'b00000000000000000000000000000000;
            code_mem[192] <= 32'b00000000000000000000000000000000;
            code_mem[193] <= 32'b00000000000000000000000000000000;
            code_mem[194] <= 32'b00000000000000000000000000000000;
            code_mem[195] <= 32'b00000000000000000000000000000000;
            code_mem[196] <= 32'b00000000000000000000000000000000;
            code_mem[197] <= 32'b00000000000000000000000000000000;
            code_mem[198] <= 32'b00000000000000000000000000000000;
            code_mem[199] <= 32'b00000000000000000000000000000000;
            code_mem[200] <= 32'b00000000000000000000000000000000;
            code_mem[201] <= 32'b00000000000000000000000000000000;
            code_mem[202] <= 32'b00000000000000000000000000000000;
            code_mem[203] <= 32'b00000000000000000000000000000000;
            code_mem[204] <= 32'b00000000000000000000000000000000;
            code_mem[205] <= 32'b00000000000000000000000000000000;
            code_mem[206] <= 32'b00000000000000000000000000000000;
            code_mem[207] <= 32'b00000000000000000000000000000000;
            code_mem[208] <= 32'b00000000000000000000000000000000;
            code_mem[209] <= 32'b00000000000000000000000000000000;
            code_mem[210] <= 32'b00000000000000000000000000000000;
            code_mem[211] <= 32'b00000000000000000000000000000000;
            code_mem[212] <= 32'b00000000000000000000000000000000;
            code_mem[213] <= 32'b00000000000000000000000000000000;
            code_mem[214] <= 32'b00000000000000000000000000000000;
            code_mem[215] <= 32'b00000000000000000000000000000000;
            code_mem[216] <= 32'b00000000000000000000000000000000;
            code_mem[217] <= 32'b00000000000000000000000000000000;
            code_mem[218] <= 32'b00000000000000000000000000000000;
            code_mem[219] <= 32'b00000000000000000000000000000000;
            code_mem[220] <= 32'b00000000000000000000000000000000;
            code_mem[221] <= 32'b00000000000000000000000000000000;
            code_mem[222] <= 32'b00000000000000000000000000000000;
            code_mem[223] <= 32'b00000000000000000000000000000000;
            code_mem[224] <= 32'b00000000000000000000000000000000;
            code_mem[225] <= 32'b00000000000000000000000000000000;
            code_mem[226] <= 32'b00000000000000000000000000000000;
            code_mem[227] <= 32'b00000000000000000000000000000000;
            code_mem[228] <= 32'b00000000000000000000000000000000;
            code_mem[229] <= 32'b00000000000000000000000000000000;
            code_mem[230] <= 32'b00000000000000000000000000000000;
            code_mem[231] <= 32'b00000000000000000000000000000000;
            code_mem[232] <= 32'b00000000000000000000000000000000;
            code_mem[233] <= 32'b00000000000000000000000000000000;
            code_mem[234] <= 32'b00000000000000000000000000000000;
            code_mem[235] <= 32'b00000000000000000000000000000000;
            code_mem[236] <= 32'b00000000000000000000000000000000;
            code_mem[237] <= 32'b00000000000000000000000000000000;
            code_mem[238] <= 32'b00000000000000000000000000000000;
            code_mem[239] <= 32'b00000000000000000000000000000000;
            code_mem[240] <= 32'b00000000000000000000000000000000;
            code_mem[241] <= 32'b00000000000000000000000000000000;
            code_mem[242] <= 32'b00000000000000000000000000000000;
            code_mem[243] <= 32'b00000000000000000000000000000000;
            code_mem[244] <= 32'b00000000000000000000000000000000;
            code_mem[245] <= 32'b00000000000000000000000000000000;
            code_mem[246] <= 32'b00000000000000000000000000000000;
            code_mem[247] <= 32'b00000000000000000000000000000000;
            code_mem[248] <= 32'b00000000000000000000000000000000;
            code_mem[249] <= 32'b00000000000000000000000000000000;
            code_mem[250] <= 32'b00000000000000000000000000000000;
            code_mem[251] <= 32'b00000000000000000000000000000000;
            code_mem[252] <= 32'b00000000000000000000000000000000;
            code_mem[253] <= 32'b00000000000000000000000000000000;
            code_mem[254] <= 32'b00000000000000000000000000000000;
            code_mem[255] <= 32'b00000000000000000000000000000000;
        end
endmodule
