`timescale 1ns / 1ps
`include "def.v"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:04:41 11/21/2018 
// Design Name: 
// Module Name:    DataMem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DataMem(
    input CLK,
    input [31:0] addr,
    input [31:0] data,
    input [5:0] opcode,
    output [31:0] out
    );
	 reg [31:0] data_mem[255:0];
	 
	 reg [31:0] read_data;
	 assign out = read_data;
	 integer i;
	 
	 always@(posedge CLK)
	  begin
			read_data <= data_mem[addr];
		end
		
	 always@(negedge CLK)
	  begin
	   if(opcode == `SDW)
			data_mem[addr] <= data;
	  end

	  initial
        begin
				read_data <= 32'b00000000000000000000000000000000;
            data_mem[0] <= 32'b00000000000000000000000000000000;
            data_mem[1] <= 32'b00000000000000000000000000000001;
            data_mem[2] <= 32'b00000000000000000000000000000010;
            data_mem[3] <= 32'b00000000000000000000000000000011;
            data_mem[4] <= 32'b00000000000000000000000000000100;
            data_mem[5] <= 32'b00000000000000000000000000000101;
            data_mem[6] <= 32'b00000000000000000000000000000110;
            data_mem[7] <= 32'b00000000000000000000000000000111;
            data_mem[8] <= 32'b00000000000000000000000000001000;
            data_mem[9] <= 32'b00000000000000000000000000001001;
            data_mem[10] <= 32'b00000000000000000000000000001010;
            data_mem[11] <= 32'b00000000000000000000000000001011;
            data_mem[12] <= 32'b00000000000000000000000000001100;
            data_mem[13] <= 32'b00000000000000000000000000001101;
            data_mem[14] <= 32'b00000000000000000000000000001110;
            data_mem[15] <= 32'b00000000000000000000000000001111;
            data_mem[16] <= 32'b00000000000000000000000000010000;
            data_mem[17] <= 32'b00000000000000000000000000010001;
            data_mem[18] <= 32'b00000000000000000000000000010010;
            data_mem[19] <= 32'b00000000000000000000000000010011;
            data_mem[20] <= 32'b00000000000000000000000000010100;
            data_mem[21] <= 32'b00000000000000000000000000010101;
            data_mem[22] <= 32'b00000000000000000000000000010110;
            data_mem[23] <= 32'b00000000000000000000000000010111;
            data_mem[24] <= 32'b00000000000000000000000000011000;
            data_mem[25] <= 32'b00000000000000000000000000011001;
            data_mem[26] <= 32'b00000000000000000000000000011010;
            data_mem[27] <= 32'b00000000000000000000000000011011;
            data_mem[28] <= 32'b00000000000000000000000000011100;
            data_mem[29] <= 32'b00000000000000000000000000011101;
            data_mem[30] <= 32'b00000000000000000000000000011110;
            data_mem[31] <= 32'b00000000000000000000000000011111;
            data_mem[32] <= 32'b00000000000000000000000000100000;
            data_mem[33] <= 32'b00000000000000000000000000100001;
            data_mem[34] <= 32'b00000000000000000000000000100010;
            data_mem[35] <= 32'b00000000000000000000000000100011;
            data_mem[36] <= 32'b00000000000000000000000000100100;
            data_mem[37] <= 32'b00000000000000000000000000100101;
            data_mem[38] <= 32'b00000000000000000000000000100110;
            data_mem[39] <= 32'b00000000000000000000000000100111;
            data_mem[40] <= 32'b00000000000000000000000000101000;
            data_mem[41] <= 32'b00000000000000000000000000101001;
            data_mem[42] <= 32'b00000000000000000000000000101010;
            data_mem[43] <= 32'b00000000000000000000000000101011;
            data_mem[44] <= 32'b00000000000000000000000000101100;
            data_mem[45] <= 32'b00000000000000000000000000101101;
            data_mem[46] <= 32'b00000000000000000000000000101110;
            data_mem[47] <= 32'b00000000000000000000000000101111;
            data_mem[48] <= 32'b00000000000000000000000000110000;
            data_mem[49] <= 32'b00000000000000000000000000110001;
            data_mem[50] <= 32'b00000000000000000000000000110010;
            data_mem[51] <= 32'b00000000000000000000000000110011;
            data_mem[52] <= 32'b00000000000000000000000000110100;
            data_mem[53] <= 32'b00000000000000000000000000110101;
            data_mem[54] <= 32'b00000000000000000000000000110110;
            data_mem[55] <= 32'b00000000000000000000000000110111;
            data_mem[56] <= 32'b00000000000000000000000000111000;
            data_mem[57] <= 32'b00000000000000000000000000111001;
            data_mem[58] <= 32'b00000000000000000000000000111010;
            data_mem[59] <= 32'b00000000000000000000000000111011;
            data_mem[60] <= 32'b00000000000000000000000000111100;
            data_mem[61] <= 32'b00000000000000000000000000111101;
            data_mem[62] <= 32'b00000000000000000000000000111110;
            data_mem[63] <= 32'b00000000000000000000000000111111;
            data_mem[64] <= 32'b00000000000000000000000001000000;
            data_mem[65] <= 32'b00000000000000000000000001000001;
            data_mem[66] <= 32'b00000000000000000000000001000010;
            data_mem[67] <= 32'b00000000000000000000000001000011;
            data_mem[68] <= 32'b00000000000000000000000001000100;
            data_mem[69] <= 32'b00000000000000000000000001000101;
            data_mem[70] <= 32'b00000000000000000000000001000110;
            data_mem[71] <= 32'b00000000000000000000000001000111;
            data_mem[72] <= 32'b00000000000000000000000001001000;
            data_mem[73] <= 32'b00000000000000000000000001001001;
            data_mem[74] <= 32'b00000000000000000000000001001010;
            data_mem[75] <= 32'b00000000000000000000000001001011;
            data_mem[76] <= 32'b00000000000000000000000001001100;
            data_mem[77] <= 32'b00000000000000000000000001001101;
            data_mem[78] <= 32'b00000000000000000000000001001110;
            data_mem[79] <= 32'b00000000000000000000000001001111;
            data_mem[80] <= 32'b00000000000000000000000001010000;
            data_mem[81] <= 32'b00000000000000000000000001010001;
            data_mem[82] <= 32'b00000000000000000000000001010010;
            data_mem[83] <= 32'b00000000000000000000000001010011;
            data_mem[84] <= 32'b00000000000000000000000001010100;
            data_mem[85] <= 32'b00000000000000000000000001010101;
            data_mem[86] <= 32'b00000000000000000000000001010110;
            data_mem[87] <= 32'b00000000000000000000000001010111;
            data_mem[88] <= 32'b00000000000000000000000001011000;
            data_mem[89] <= 32'b00000000000000000000000001011001;
            data_mem[90] <= 32'b00000000000000000000000001011010;
            data_mem[91] <= 32'b00000000000000000000000001011011;
            data_mem[92] <= 32'b00000000000000000000000001011100;
            data_mem[93] <= 32'b00000000000000000000000001011101;
            data_mem[94] <= 32'b00000000000000000000000001011110;
            data_mem[95] <= 32'b00000000000000000000000001011111;
            data_mem[96] <= 32'b00000000000000000000000001100000;
            data_mem[97] <= 32'b00000000000000000000000001100001;
            data_mem[98] <= 32'b00000000000000000000000001100010;
            data_mem[99] <= 32'b00000000000000000000000001100011;
            data_mem[100] <= 32'b00000000000000000000000001100100;
            data_mem[101] <= 32'b00000000000000000000000001100101;
            data_mem[102] <= 32'b00000000000000000000000001100110;
            data_mem[103] <= 32'b00000000000000000000000001100111;
            data_mem[104] <= 32'b00000000000000000000000001101000;
            data_mem[105] <= 32'b00000000000000000000000001101001;
            data_mem[106] <= 32'b00000000000000000000000001101010;
            data_mem[107] <= 32'b00000000000000000000000001101011;
            data_mem[108] <= 32'b00000000000000000000000001101100;
            data_mem[109] <= 32'b00000000000000000000000001101101;
            data_mem[110] <= 32'b00000000000000000000000001101110;
            data_mem[111] <= 32'b00000000000000000000000001101111;
            data_mem[112] <= 32'b00000000000000000000000001110000;
            data_mem[113] <= 32'b00000000000000000000000001110001;
            data_mem[114] <= 32'b00000000000000000000000001110010;
            data_mem[115] <= 32'b00000000000000000000000001110011;
            data_mem[116] <= 32'b00000000000000000000000001110100;
            data_mem[117] <= 32'b00000000000000000000000001110101;
            data_mem[118] <= 32'b00000000000000000000000001110110;
            data_mem[119] <= 32'b00000000000000000000000001110111;
            data_mem[120] <= 32'b00000000000000000000000001111000;
            data_mem[121] <= 32'b00000000000000000000000001111001;
            data_mem[122] <= 32'b00000000000000000000000001111010;
            data_mem[123] <= 32'b00000000000000000000000001111011;
            data_mem[124] <= 32'b00000000000000000000000001111100;
            data_mem[125] <= 32'b00000000000000000000000001111101;
            data_mem[126] <= 32'b00000000000000000000000001111110;
            data_mem[127] <= 32'b00000000000000000000000001111111;
            data_mem[128] <= 32'b00000000000000000000000010000000;
            data_mem[129] <= 32'b00000000000000000000000010000001;
            data_mem[130] <= 32'b00000000000000000000000010000010;
            data_mem[131] <= 32'b00000000000000000000000010000011;
            data_mem[132] <= 32'b00000000000000000000000010000100;
            data_mem[133] <= 32'b00000000000000000000000010000101;
            data_mem[134] <= 32'b00000000000000000000000010000110;
            data_mem[135] <= 32'b00000000000000000000000010000111;
            data_mem[136] <= 32'b00000000000000000000000010001000;
            data_mem[137] <= 32'b00000000000000000000000010001001;
            data_mem[138] <= 32'b00000000000000000000000010001010;
            data_mem[139] <= 32'b00000000000000000000000010001011;
            data_mem[140] <= 32'b00000000000000000000000010001100;
            data_mem[141] <= 32'b00000000000000000000000010001101;
            data_mem[142] <= 32'b00000000000000000000000010001110;
            data_mem[143] <= 32'b00000000000000000000000010001111;
            data_mem[144] <= 32'b00000000000000000000000010010000;
            data_mem[145] <= 32'b00000000000000000000000010010001;
            data_mem[146] <= 32'b00000000000000000000000010010010;
            data_mem[147] <= 32'b00000000000000000000000010010011;
            data_mem[148] <= 32'b00000000000000000000000010010100;
            data_mem[149] <= 32'b00000000000000000000000010010101;
            data_mem[150] <= 32'b00000000000000000000000010010110;
            data_mem[151] <= 32'b00000000000000000000000010010111;
            data_mem[152] <= 32'b00000000000000000000000010011000;
            data_mem[153] <= 32'b00000000000000000000000010011001;
            data_mem[154] <= 32'b00000000000000000000000010011010;
            data_mem[155] <= 32'b00000000000000000000000010011011;
            data_mem[156] <= 32'b00000000000000000000000010011100;
            data_mem[157] <= 32'b00000000000000000000000010011101;
            data_mem[158] <= 32'b00000000000000000000000010011110;
            data_mem[159] <= 32'b00000000000000000000000010011111;
            data_mem[160] <= 32'b00000000000000000000000010100000;
            data_mem[161] <= 32'b00000000000000000000000010100001;
            data_mem[162] <= 32'b00000000000000000000000010100010;
            data_mem[163] <= 32'b00000000000000000000000010100011;
            data_mem[164] <= 32'b00000000000000000000000010100100;
            data_mem[165] <= 32'b00000000000000000000000010100101;
            data_mem[166] <= 32'b00000000000000000000000010100110;
            data_mem[167] <= 32'b00000000000000000000000010100111;
            data_mem[168] <= 32'b00000000000000000000000010101000;
            data_mem[169] <= 32'b00000000000000000000000010101001;
            data_mem[170] <= 32'b00000000000000000000000010101010;
            data_mem[171] <= 32'b00000000000000000000000010101011;
            data_mem[172] <= 32'b00000000000000000000000010101100;
            data_mem[173] <= 32'b00000000000000000000000010101101;
            data_mem[174] <= 32'b00000000000000000000000010101110;
            data_mem[175] <= 32'b00000000000000000000000010101111;
            data_mem[176] <= 32'b00000000000000000000000010110000;
            data_mem[177] <= 32'b00000000000000000000000010110001;
            data_mem[178] <= 32'b00000000000000000000000010110010;
            data_mem[179] <= 32'b00000000000000000000000010110011;
            data_mem[180] <= 32'b00000000000000000000000010110100;
            data_mem[181] <= 32'b00000000000000000000000010110101;
            data_mem[182] <= 32'b00000000000000000000000010110110;
            data_mem[183] <= 32'b00000000000000000000000010110111;
            data_mem[184] <= 32'b00000000000000000000000010111000;
            data_mem[185] <= 32'b00000000000000000000000010111001;
            data_mem[186] <= 32'b00000000000000000000000010111010;
            data_mem[187] <= 32'b00000000000000000000000010111011;
            data_mem[188] <= 32'b00000000000000000000000010111100;
            data_mem[189] <= 32'b00000000000000000000000010111101;
            data_mem[190] <= 32'b00000000000000000000000010111110;
            data_mem[191] <= 32'b00000000000000000000000010111111;
            data_mem[192] <= 32'b00000000000000000000000011000000;
            data_mem[193] <= 32'b00000000000000000000000011000001;
            data_mem[194] <= 32'b00000000000000000000000011000010;
            data_mem[195] <= 32'b00000000000000000000000011000011;
            data_mem[196] <= 32'b00000000000000000000000011000100;
            data_mem[197] <= 32'b00000000000000000000000011000101;
            data_mem[198] <= 32'b00000000000000000000000011000110;
            data_mem[199] <= 32'b00000000000000000000000011000111;
            data_mem[200] <= 32'b00000000000000000000000011001000;
            data_mem[201] <= 32'b00000000000000000000000011001001;
            data_mem[202] <= 32'b00000000000000000000000011001010;
            data_mem[203] <= 32'b00000000000000000000000011001011;
            data_mem[204] <= 32'b00000000000000000000000011001100;
            data_mem[205] <= 32'b00000000000000000000000011001101;
            data_mem[206] <= 32'b00000000000000000000000011001110;
            data_mem[207] <= 32'b00000000000000000000000011001111;
            data_mem[208] <= 32'b00000000000000000000000011010000;
            data_mem[209] <= 32'b00000000000000000000000011010001;
            data_mem[210] <= 32'b00000000000000000000000011010010;
            data_mem[211] <= 32'b00000000000000000000000011010011;
            data_mem[212] <= 32'b00000000000000000000000011010100;
            data_mem[213] <= 32'b00000000000000000000000011010101;
            data_mem[214] <= 32'b00000000000000000000000011010110;
            data_mem[215] <= 32'b00000000000000000000000011010111;
            data_mem[216] <= 32'b00000000000000000000000011011000;
            data_mem[217] <= 32'b00000000000000000000000011011001;
            data_mem[218] <= 32'b00000000000000000000000011011010;
            data_mem[219] <= 32'b00000000000000000000000011011011;
            data_mem[220] <= 32'b00000000000000000000000011011100;
            data_mem[221] <= 32'b00000000000000000000000011011101;
            data_mem[222] <= 32'b00000000000000000000000011011110;
            data_mem[223] <= 32'b00000000000000000000000011011111;
            data_mem[224] <= 32'b00000000000000000000000011100000;
            data_mem[225] <= 32'b00000000000000000000000011100001;
            data_mem[226] <= 32'b00000000000000000000000011100010;
            data_mem[227] <= 32'b00000000000000000000000011100011;
            data_mem[228] <= 32'b00000000000000000000000011100100;
            data_mem[229] <= 32'b00000000000000000000000011100101;
            data_mem[230] <= 32'b00000000000000000000000011100110;
            data_mem[231] <= 32'b00000000000000000000000011100111;
            data_mem[232] <= 32'b00000000000000000000000011101000;
            data_mem[233] <= 32'b00000000000000000000000011101001;
            data_mem[234] <= 32'b00000000000000000000000011101010;
            data_mem[235] <= 32'b00000000000000000000000011101011;
            data_mem[236] <= 32'b00000000000000000000000011101100;
            data_mem[237] <= 32'b00000000000000000000000011101101;
            data_mem[238] <= 32'b00000000000000000000000011101110;
            data_mem[239] <= 32'b00000000000000000000000011101111;
            data_mem[240] <= 32'b00000000000000000000000011110000;
            data_mem[241] <= 32'b00000000000000000000000011110001;
            data_mem[242] <= 32'b00000000000000000000000011110010;
            data_mem[243] <= 32'b00000000000000000000000011110011;
            data_mem[244] <= 32'b00000000000000000000000011110100;
            data_mem[245] <= 32'b00000000000000000000000011110101;
            data_mem[246] <= 32'b00000000000000000000000011110110;
            data_mem[247] <= 32'b00000000000000000000000011110111;
            data_mem[248] <= 32'b00000000000000000000000011111000;
            data_mem[249] <= 32'b00000000000000000000000011111001;
            data_mem[250] <= 32'b00000000000000000000000011111010;
            data_mem[251] <= 32'b00000000000000000000000011111011;
            data_mem[252] <= 32'b00000000000000000000000011111100;
            data_mem[253] <= 32'b00000000000000000000000011111101;
            data_mem[254] <= 32'b00000000000000000000000011111110;
				data_mem[255] <= 32'b00000000000000000000000011111111;
        end
endmodule
